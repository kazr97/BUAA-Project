`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:55:33 12/10/2017 
// Design Name: 
// Module Name:    control 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
	module control(
	input [31:0] IR,
	input [5:0] op,func,
	output reg EXTsle,MUX_ALU_B_sle,RegWrite,Branch,ifj,start,M,cp,eret,WA,
	output reg [1:0] MUX_A3_sle,MUX_WDOUT_sle,npcsle,MemWrite,
	output reg [2:0] CMPsle,
	output reg [3:0] ALUsle,kuo,MULTsle
    );
	always @ *begin
		case(op)
			6'b000000:begin
				case(func)
					6'b100001:begin
						EXTsle<=0;
						npcsle<=0;
						MUX_ALU_B_sle<=0;
						ALUsle<=0;
						RegWrite<=1;
						Branch<=0;
						MUX_A3_sle<=1;
						MUX_WDOUT_sle<=0;
						MemWrite<=0;
						CMPsle<=0;
						ifj<=0;
						kuo<=0;
						start<=0;
						MULTsle<=0;
						M<=0;
						cp<=0;
						eret<=0;
						WA<=0;
					end//addu
					
					6'b100000:begin
						EXTsle<=0;
						npcsle<=0;
						MUX_ALU_B_sle<=0;
						ALUsle<=0;
						RegWrite<=1;
						Branch<=0;
						MUX_A3_sle<=1;
						MUX_WDOUT_sle<=0;
						MemWrite<=0;
						CMPsle<=0;
						ifj<=0;
						kuo<=0;
						start<=0;
						MULTsle<=0;
						M<=0;
						cp<=0;
						eret<=0;
						WA<=0;
					end//add
					
					6'b100011:begin
						EXTsle<=0;
						npcsle<=0;
						MUX_ALU_B_sle<=0;
						ALUsle<=1;
						RegWrite<=1;
						Branch<=0;
						MUX_A3_sle<=1;
						MUX_WDOUT_sle<=0;
						MemWrite<=0;
						CMPsle<=0;
						ifj<=0;
						kuo<=0;
						start<=0;
						MULTsle<=0;
						M<=0;
						cp<=0;
						eret<=0;
						WA<=0;
					end//subu
					
					6'b100010:begin
						EXTsle<=0;
						npcsle<=0;
						MUX_ALU_B_sle<=0;
						ALUsle<=1;
						RegWrite<=1;
						Branch<=0;
						MUX_A3_sle<=1;
						MUX_WDOUT_sle<=0;
						MemWrite<=0;
						CMPsle<=0;
						ifj<=0;
						kuo<=0;
						start<=0;
						MULTsle<=0;
						M<=0;
						cp<=0;
						eret<=0;
						WA<=0;
					end//sub
					
					6'b001000:begin
						EXTsle<=0;
						npcsle<=3;
						MUX_ALU_B_sle<=0;
						ALUsle<=0;
						RegWrite<=0;
						Branch<=0;
						MUX_A3_sle<=0;
						MUX_WDOUT_sle<=0;
						MemWrite<=0;
						CMPsle<=0;
						ifj<=1;
						kuo<=0;
						start<=0;
						MULTsle<=0;
						M<=0;
						cp<=0;
						eret<=0;
						WA<=0;
					end//jr
					
					6'b001001:begin
						EXTsle<=0;
						npcsle<=3;
						MUX_ALU_B_sle<=0;
						ALUsle<=4;
						RegWrite<=1;
						Branch<=0;
						MUX_A3_sle<=1;
						MUX_WDOUT_sle<=2;
						MemWrite<=0;
						CMPsle<=0;
						ifj<=1;
						kuo<=0;
						start<=0;
						MULTsle<=0;
						M<=0;
						cp<=0;
						eret<=0;
						WA<=0;
					end//jalr
					
					6'b000000:begin
						EXTsle<=0;
						npcsle<=0;
						MUX_ALU_B_sle<=0;
						ALUsle<=5;
						RegWrite<=1;
						Branch<=0;
						MUX_A3_sle<=1;
						MUX_WDOUT_sle<=0;
						MemWrite<=0;
						CMPsle<=0;
						ifj<=0;
						kuo<=0;
						start<=0;
						MULTsle<=0;
						M<=0;
						cp<=0;
						eret<=0;
						WA<=0;
					end//sll
					
					6'b000010:begin
						EXTsle<=0;
						npcsle<=0;
						MUX_ALU_B_sle<=0;
						ALUsle<=6;
						RegWrite<=1;
						Branch<=0;
						MUX_A3_sle<=1;
						MUX_WDOUT_sle<=0;
						MemWrite<=0;
						CMPsle<=0;
						ifj<=0;
						kuo<=0;
						start<=0;
						MULTsle<=0;
						M<=0;
						cp<=0;
						eret<=0;
						WA<=0;
					end//srl
					
					6'b000011:begin
						EXTsle<=0;
						npcsle<=0;
						MUX_ALU_B_sle<=0;
						ALUsle<=7;
						RegWrite<=1;
						Branch<=0;
						MUX_A3_sle<=1;
						MUX_WDOUT_sle<=0;
						MemWrite<=0;
						CMPsle<=0;
						ifj<=0;
						kuo<=0;
						start<=0;
						MULTsle<=0;
						M<=0;
						cp<=0;
						eret<=0;
						WA<=0;
					end//sra
					
					6'b000100:begin
						EXTsle<=0;
						npcsle<=0;
						MUX_ALU_B_sle<=0;
						ALUsle<=8;
						RegWrite<=1;
						Branch<=0;
						MUX_A3_sle<=1;
						MUX_WDOUT_sle<=0;
						MemWrite<=0;
						CMPsle<=0;
						ifj<=0;
						kuo<=0;
						start<=0;
						MULTsle<=0;
						M<=0;
						cp<=0;
						eret<=0;
						WA<=0;
					end//sllv
					
					6'b000110:begin
						EXTsle<=0;
						npcsle<=0;
						MUX_ALU_B_sle<=0;
						ALUsle<=9;
						RegWrite<=1;
						Branch<=0;
						MUX_A3_sle<=1;
						MUX_WDOUT_sle<=0;
						MemWrite<=0;
						CMPsle<=0;
						ifj<=0;
						kuo<=0;
						start<=0;
						MULTsle<=0;
						M<=0;
						cp<=0;
						eret<=0;
						WA<=0;
					end//srlv
					
					6'b000111:begin
						EXTsle<=0;
						npcsle<=0;
						MUX_ALU_B_sle<=0;
						ALUsle<=10;
						RegWrite<=1;
						Branch<=0;
						MUX_A3_sle<=1;
						MUX_WDOUT_sle<=0;
						MemWrite<=0;
						CMPsle<=0;
						ifj<=0;
						kuo<=0;
						start<=0;
						MULTsle<=0;
						M<=0;
						cp<=0;
						eret<=0;
						WA<=0;
					end//srav
					
					6'b100100:begin
						EXTsle<=1;
						npcsle<=0;
						MUX_ALU_B_sle<=0;
						ALUsle<=11;
						RegWrite<=1;
						Branch<=0;
						MUX_A3_sle<=1;
						MUX_WDOUT_sle<=0;
						MemWrite<=0;
						CMPsle<=0;
						ifj<=0;
						kuo<=0;
						start<=0;
						MULTsle<=0;
						M<=0;
						cp<=0;
						eret<=0;
						WA<=0;
					end//and
					
					6'b100101:begin
						EXTsle<=1;
						npcsle<=0;
						MUX_ALU_B_sle<=0;
						ALUsle<=2;
						RegWrite<=1;
						Branch<=0;
						MUX_A3_sle<=1;
						MUX_WDOUT_sle<=0;
						MemWrite<=0;
						CMPsle<=0;
						ifj<=0;
						kuo<=0;
						start<=0;
						MULTsle<=0;
						M<=0;
						cp<=0;
						eret<=0;
						WA<=0;
					end//or
					
					6'b100110:begin
						EXTsle<=1;
						npcsle<=0;
						MUX_ALU_B_sle<=0;
						ALUsle<=12;
						RegWrite<=1;
						Branch<=0;
						MUX_A3_sle<=1;
						MUX_WDOUT_sle<=0;
						MemWrite<=0;
						CMPsle<=0;
						ifj<=0;
						kuo<=0;
						start<=0;
						MULTsle<=0;
						M<=0;
						cp<=0;
						eret<=0;
						WA<=0;
					end//xor
					
					6'b100111:begin
						EXTsle<=1;
						npcsle<=0;
						MUX_ALU_B_sle<=0;
						ALUsle<=13;
						RegWrite<=1;
						Branch<=0;
						MUX_A3_sle<=1;
						MUX_WDOUT_sle<=0;
						MemWrite<=0;
						CMPsle<=0;
						ifj<=0;
						kuo<=0;
						start<=0;
						MULTsle<=0;
						M<=0;
						cp<=0;
						eret<=0;
						WA<=0;
					end//nor
					
					6'b101010:begin
						EXTsle<=0;
						npcsle<=0;
						MUX_ALU_B_sle<=0;
						ALUsle<=14;
						RegWrite<=1;
						Branch<=0;
						MUX_A3_sle<=1;
						MUX_WDOUT_sle<=0;
						MemWrite<=0;
						CMPsle<=0;
						ifj<=0;
						kuo<=0;
						start<=0;
						MULTsle<=0;
						M<=0;
						cp<=0;
						eret<=0;
						WA<=0;
					end//slt
					
					6'b101011:begin
						EXTsle<=0;
						npcsle<=0;
						MUX_ALU_B_sle<=0;
						ALUsle<=15;
						RegWrite<=1;
						Branch<=0;
						MUX_A3_sle<=1;
						MUX_WDOUT_sle<=0;
						MemWrite<=0;
						CMPsle<=0;
						ifj<=0;
						kuo<=0;
						start<=0;
						MULTsle<=0;
						M<=0;
						cp<=0;
						eret<=0;
						WA<=0;
					end//sltu
					
					6'b011000:begin
						EXTsle<=0;
						npcsle<=0;
						MUX_ALU_B_sle<=0;
						ALUsle<=0;
						RegWrite<=0;
						Branch<=0;
						MUX_A3_sle<=0;
						MUX_WDOUT_sle<=0;
						MemWrite<=0;
						CMPsle<=0;
						ifj<=0;
						kuo<=0;
						start<=1;
						MULTsle<=0;
						M<=1;
						cp<=0;
						eret<=0;
						WA<=0;
					end//mult
					
					6'b011001:begin
						EXTsle<=0;
						npcsle<=0;
						MUX_ALU_B_sle<=0;
						ALUsle<=0;
						RegWrite<=0;
						Branch<=0;
						MUX_A3_sle<=0;
						MUX_WDOUT_sle<=0;
						MemWrite<=0;
						CMPsle<=0;
						ifj<=0;
						kuo<=0;
						start<=1;
						MULTsle<=1;
						M<=1;
						cp<=0;
						eret<=0;
						WA<=0;
					end//multu
					
					6'b011010:begin
						EXTsle<=0;
						npcsle<=0;
						MUX_ALU_B_sle<=0;
						ALUsle<=0;
						RegWrite<=0;
						Branch<=0;
						MUX_A3_sle<=0;
						MUX_WDOUT_sle<=0;
						MemWrite<=0;
						CMPsle<=0;
						ifj<=0;
						kuo<=0;
						start<=1;
						MULTsle<=2;
						M<=1;
						cp<=0;
						eret<=0;
						WA<=0;
					end//div
					
					6'b011011:begin
						EXTsle<=0;
						npcsle<=0;
						MUX_ALU_B_sle<=0;
						ALUsle<=0;
						RegWrite<=0;
						Branch<=0;
						MUX_A3_sle<=0;
						MUX_WDOUT_sle<=0;
						MemWrite<=0;
						CMPsle<=0;
						ifj<=0;
						kuo<=0;
						start<=1;
						MULTsle<=3;
						M<=1;
						cp<=0;
						eret<=0;
						WA<=0;
					end//divu
					
					6'b010000:begin
						EXTsle<=0;
						npcsle<=0;
						MUX_ALU_B_sle<=0;
						ALUsle<=0;
						RegWrite<=1;
						Branch<=0;
						MUX_A3_sle<=1;
						MUX_WDOUT_sle<=0;
						MemWrite<=0;
						CMPsle<=0;
						ifj<=0;
						kuo<=0;
						start<=0;
						MULTsle<=4;
						M<=1;
						cp<=0;
						eret<=0;
						WA<=0;
					end//mfhi
					
					6'b010010:begin
						EXTsle<=0;
						npcsle<=0;
						MUX_ALU_B_sle<=0;
						ALUsle<=0;
						RegWrite<=1;
						Branch<=0;
						MUX_A3_sle<=1;
						MUX_WDOUT_sle<=0;
						MemWrite<=0;
						CMPsle<=0;
						ifj<=0;
						kuo<=0;
						start<=0;
						MULTsle<=5;
						M<=1;
						cp<=0;
						eret<=0;
						WA<=0;
					end//mflo
					
					6'b010001:begin
						EXTsle<=0;
						npcsle<=0;
						MUX_ALU_B_sle<=0;
						ALUsle<=0;
						RegWrite<=0;
						Branch<=0;
						MUX_A3_sle<=0;
						MUX_WDOUT_sle<=0;
						MemWrite<=0;
						CMPsle<=0;
						ifj<=0;
						kuo<=0;
						start<=0;
						MULTsle<=6;
						M<=1;
						cp<=0;
						eret<=0;
						WA<=0;
					end//mthi
					
					6'b010011:begin
						EXTsle<=0;
						npcsle<=0;
						MUX_ALU_B_sle<=0;
						ALUsle<=0;
						RegWrite<=0;
						Branch<=0;
						MUX_A3_sle<=0;
						MUX_WDOUT_sle<=0;
						MemWrite<=0;
						CMPsle<=0;
						ifj<=0;
						kuo<=0;
						start<=0;
						MULTsle<=7;
						M<=1;
						cp<=0;
						eret<=0;
						WA<=0;
					end//mthi
					
					6'b000000:begin
						EXTsle<=0;
						npcsle<=0;
						MUX_ALU_B_sle<=0;
						ALUsle<=0;
						RegWrite<=0;
						Branch<=0;
						MUX_A3_sle<=0;
						MUX_WDOUT_sle<=0;
						MemWrite<=0;
						CMPsle<=0;
						ifj<=0;
						kuo<=0;
						start<=0;
						MULTsle<=0;
						M<=0;
						cp<=0;
						eret<=0;
						WA<=0;
					end//nop

					
					default begin
						EXTsle<=0;
						npcsle<=0;
						MUX_ALU_B_sle<=0;
						ALUsle<=0;
						RegWrite<=0;
						Branch<=0;
						MUX_A3_sle<=0;
						MUX_WDOUT_sle<=0;
						MemWrite<=0;
						CMPsle<=0;
						ifj<=0;
						kuo<=0;
						start<=0;
						MULTsle<=0;
						M<=0;
						cp<=0;
						eret<=0;
						WA<=1;
					end
				endcase
			end
			
			6'b001101:begin
				EXTsle<=1;
				npcsle<=0;
				MUX_ALU_B_sle<=1;
				ALUsle<=2;
				RegWrite<=1;
				Branch<=0;
				MUX_A3_sle<=0;
				MUX_WDOUT_sle<=0;
				MemWrite<=0;
				CMPsle<=0;
				ifj<=0;
				kuo<=0;
				start<=0;
				MULTsle<=0;
				M<=0;
				cp<=0;
				eret<=0;
				WA<=0;
			end//ori
			
			6'b100011:begin
				EXTsle<=0;
				npcsle<=0;
				MUX_ALU_B_sle<=1;
				ALUsle<=0;
				RegWrite<=1;
				Branch<=0;
				MUX_A3_sle<=0;
				MUX_WDOUT_sle<=1;
				MemWrite<=0;
				CMPsle<=0;
				ifj<=0;
				kuo<=0;
				start<=0;
				MULTsle<=0;
				M<=0;
				cp<=0;
				eret<=0;
				WA<=0;
			end//lw
			
			6'b101011:begin
				EXTsle<=0;
				npcsle<=0;
				MUX_ALU_B_sle<=1;
				ALUsle<=0;
				RegWrite<=0;
				Branch<=0;
				MUX_A3_sle<=0;
				MUX_WDOUT_sle<=0;
				MemWrite<=1;
				CMPsle<=0;
				ifj<=0;
				kuo<=0;
				start<=0;
				MULTsle<=0;
				M<=0;
				cp<=0;
				eret<=0;
				WA<=0;
			end//sw
			
			6'b000100:begin
				EXTsle<=0;
				npcsle<=1;
				MUX_ALU_B_sle<=0;
				ALUsle<=0;
				RegWrite<=0;
				Branch<=1;
				MUX_A3_sle<=0;
				MUX_WDOUT_sle<=0;
				MemWrite<=0;
				CMPsle<=0;
				ifj<=0;
				kuo<=0;
				start<=0;
				MULTsle<=0;
				M<=0;
				cp<=0;
				eret<=0;
				WA<=0;
			end//beq
			
			6'b001111:begin
				EXTsle<=0;
				npcsle<=0;
				MUX_ALU_B_sle<=1;
				ALUsle<=3;
				RegWrite<=1;
				Branch<=0;
				MUX_A3_sle<=0;
				MUX_WDOUT_sle<=0;
				MemWrite<=0;
				CMPsle<=0;
				ifj<=0;
				kuo<=0;
				start<=0;
				MULTsle<=0;
				M<=0;
				cp<=0;
				eret<=0;
				WA<=0;
			end//lui
			
			6'b000010:begin
				EXTsle<=0;
				npcsle<=2;
				MUX_ALU_B_sle<=1;
				ALUsle<=0;
				RegWrite<=0;
				Branch<=0;
				MUX_A3_sle<=0;
				MUX_WDOUT_sle<=0;
				MemWrite<=0;
				CMPsle<=0;
				ifj<=1;
				kuo<=0;
				start<=0;
				MULTsle<=0;
				M<=0;
				cp<=0;
				eret<=0;
				WA<=0;
			end//j
			
			6'b000011:begin
				EXTsle<=0;
				npcsle<=2;
				MUX_ALU_B_sle<=0;
				ALUsle<=4;
				RegWrite<=1;
				Branch<=0;
				MUX_A3_sle<=2;
				MUX_WDOUT_sle<=2;
				MemWrite<=0;
				CMPsle<=0;
				ifj<=1;
				kuo<=0;
				start<=0;
				MULTsle<=0;
				M<=0;
				cp<=0;
				eret<=0;
				WA<=0;
			end//jal
			
			6'b000101:begin
				EXTsle<=0;
				npcsle<=1;
				MUX_ALU_B_sle<=0;
				ALUsle<=0;
				RegWrite<=0;
				Branch<=1;
				MUX_A3_sle<=0;
				MUX_WDOUT_sle<=0;
				MemWrite<=0;
				CMPsle<=1;
				ifj<=0;
				kuo<=0;
				start<=0;
				MULTsle<=0;
				M<=0;
				cp<=0;
				eret<=0;
				WA<=0;
			end//bne
			
			6'b101001:begin
				EXTsle<=0;
				npcsle<=0;
				MUX_ALU_B_sle<=1;
				ALUsle<=0;
				RegWrite<=0;
				Branch<=0;
				MUX_A3_sle<=0;
				MUX_WDOUT_sle<=0;
				MemWrite<=2;
				CMPsle<=0;
				ifj<=0;
				kuo<=0;
				start<=0;
				MULTsle<=0;
				M<=0;
				cp<=0;
				eret<=0;
				WA<=0;
			end//////sh
				
			6'b100000:begin
				EXTsle<=0;
				npcsle<=0;
				MUX_ALU_B_sle<=1;
				ALUsle<=0;
				RegWrite<=1;
				Branch<=0;
				MUX_A3_sle<=0;
				MUX_WDOUT_sle<=1;
				MemWrite<=0;
				CMPsle<=0;
				ifj<=0;
				kuo<=4;
				start<=0;
				MULTsle<=0;
				M<=0;
				cp<=0;
				eret<=0;
				WA<=0;
			end////lb
			
			6'b100100:begin
				EXTsle<=0;
				npcsle<=0;
				MUX_ALU_B_sle<=1;
				ALUsle<=0;
				RegWrite<=1;
				Branch<=0;
				MUX_A3_sle<=0;
				MUX_WDOUT_sle<=1;
				MemWrite<=0;
				CMPsle<=0;
				ifj<=0;
				kuo<=3;
				start<=0;
				MULTsle<=0;
				M<=0;
				cp<=0;
				eret<=0;
				WA<=0;
			end/////lbu
			
			6'b100001:begin
				EXTsle<=0;
				npcsle<=0;
				MUX_ALU_B_sle<=1;
				ALUsle<=0;
				RegWrite<=1;
				Branch<=0;
				MUX_A3_sle<=0;
				MUX_WDOUT_sle<=1;
				MemWrite<=0;
				CMPsle<=0;
				ifj<=0;
				kuo<=2;
				start<=0;
				MULTsle<=0;
				M<=0;
				cp<=0;
				eret<=0;
				WA<=0;
			end/////lh
			
			6'b100101:begin
				EXTsle<=0;
				npcsle<=0;
				MUX_ALU_B_sle<=1;
				ALUsle<=0;
				RegWrite<=1;
				Branch<=0;
				MUX_A3_sle<=0;
				MUX_WDOUT_sle<=1;
				MemWrite<=0;
				CMPsle<=0;
				ifj<=0;
				kuo<=1;
				start<=0;
				MULTsle<=0;
				M<=0;
				cp<=0;
				eret<=0;
				WA<=0;
			end/////lhu
			
			6'b101000:begin
				EXTsle<=0;
				npcsle<=0;
				MUX_ALU_B_sle<=1;
				ALUsle<=0;
				RegWrite<=0;
				Branch<=0;
				MUX_A3_sle<=0;
				MUX_WDOUT_sle<=0;
				MemWrite<=3;
				CMPsle<=0;
				ifj<=0;
				kuo<=0;
				start<=0;
				MULTsle<=0;
				M<=0;
				cp<=0;
				eret<=0;
				WA<=0;
			end//////sb
			
			6'b001000:begin
				EXTsle<=0;
				npcsle<=0;
				MUX_ALU_B_sle<=1;
				ALUsle<=0;
				RegWrite<=1;
				Branch<=0;
				MUX_A3_sle<=0;
				MUX_WDOUT_sle<=0;
				MemWrite<=0;
				CMPsle<=0;
				ifj<=0;
				kuo<=0;
				start<=0;
				MULTsle<=0;
				M<=0;
				cp<=0;
				eret<=0;
				WA<=0;
			end//////addi
					
			6'b001001:begin
				EXTsle<=0;
				npcsle<=0;
				MUX_ALU_B_sle<=1;
				ALUsle<=0;
				RegWrite<=1;
				Branch<=0;
				MUX_A3_sle<=0;
				MUX_WDOUT_sle<=0;
				MemWrite<=0;
				CMPsle<=0;
				ifj<=0;
				kuo<=0;
				start<=0;
				MULTsle<=0;
				M<=0;
				cp<=0;
				eret<=0;
				WA<=0;
			end//////addiu

			6'b001100:begin
				EXTsle<=1;
				npcsle<=0;
				MUX_ALU_B_sle<=1;
				ALUsle<=11;
				RegWrite<=1;
				Branch<=0;
				MUX_A3_sle<=0;
				MUX_WDOUT_sle<=0;
				MemWrite<=0;
				CMPsle<=0;
				ifj<=0;
				kuo<=0;
				start<=0;
				MULTsle<=0;
				M<=0;
				cp<=0;
				eret<=0;
				WA<=0;
			end//////andi		

			6'b001110:begin
				EXTsle<=1;
				npcsle<=0;
				MUX_ALU_B_sle<=1;
				ALUsle<=12;
				RegWrite<=1;
				Branch<=0;
				MUX_A3_sle<=0;
				MUX_WDOUT_sle<=0;
				MemWrite<=0;
				CMPsle<=0;
				ifj<=0;
				kuo<=0;
				start<=0;
				MULTsle<=0;
				M<=0;
				cp<=0;
				eret<=0;
				WA<=0;
			end//////xori

			6'b001010:begin
				EXTsle<=0;
				npcsle<=0;
				MUX_ALU_B_sle<=1;
				ALUsle<=14;
				RegWrite<=1;
				Branch<=0;
				MUX_A3_sle<=0;
				MUX_WDOUT_sle<=0;
				MemWrite<=0;
				CMPsle<=0;
				ifj<=0;
				kuo<=0;
				start<=0;
				MULTsle<=0;
				M<=0;
				cp<=0;
				eret<=0;
				WA<=0;
			end//////slti	

			6'b001011:begin
				EXTsle<=0;
				npcsle<=0;
				MUX_ALU_B_sle<=1;
				ALUsle<=15;
				RegWrite<=1;
				Branch<=0;
				MUX_A3_sle<=0;
				MUX_WDOUT_sle<=0;
				MemWrite<=0;
				CMPsle<=0;
				ifj<=0;
				kuo<=0;
				start<=0;
				MULTsle<=0;
				M<=0;
				cp<=0;
				eret<=0;
				WA<=0;
			end//////sltiu
			
			6'b000110:begin
				EXTsle<=0;
				npcsle<=1;
				MUX_ALU_B_sle<=0;
				ALUsle<=0;
				RegWrite<=0;
				Branch<=1;
				MUX_A3_sle<=0;
				MUX_WDOUT_sle<=0;
				MemWrite<=0;
				CMPsle<=3;
				ifj<=0;
				kuo<=0;
				start<=0;
				MULTsle<=0;
				M<=0;
				cp<=0;
				eret<=0;
				WA<=0;
			end//////blez
			
			6'b000111:begin
				EXTsle<=0;
				npcsle<=1;
				MUX_ALU_B_sle<=0;
				ALUsle<=0;
				RegWrite<=0;
				Branch<=1;
				MUX_A3_sle<=0;
				MUX_WDOUT_sle<=0;
				MemWrite<=0;
				CMPsle<=4;
				ifj<=0;
				kuo<=0;
				start<=0;
				MULTsle<=0;
				M<=0;
				cp<=0;
				eret<=0;
				WA<=0;
			end//////bgtz
			
			6'b010000:begin
				case(IR[25:21])
					5'b00100:begin
						EXTsle<=0;
						npcsle<=0;
						MUX_ALU_B_sle<=0;
						ALUsle<=0;
						RegWrite<=0;
						Branch<=0;
						MUX_A3_sle<=0;
						MUX_WDOUT_sle<=0;
						MemWrite<=0;
						CMPsle<=0;
						ifj<=0;
						kuo<=0;
						start<=0;
						MULTsle<=0;
						M<=0;
						cp<=1;
						eret<=0;
						WA<=0;
					end//////mtc0
					
					5'b00000:begin
						EXTsle<=0;
						npcsle<=0;
						MUX_ALU_B_sle<=0;
						ALUsle<=0;
						RegWrite<=1;
						Branch<=0;
						MUX_A3_sle<=0;
						MUX_WDOUT_sle<=1;
						MemWrite<=0;
						CMPsle<=0;
						ifj<=0;
						kuo<=0;
						start<=0;
						MULTsle<=0;
						M<=0;
						cp<=1;
						eret<=0;
						WA<=0;
					end//////mfc0
				endcase
				
				case(func)
					6'b011000:begin
						EXTsle<=0;
						npcsle<=0;
						MUX_ALU_B_sle<=0;
						ALUsle<=0;
						RegWrite<=0;
						Branch<=0;
						MUX_A3_sle<=0;
						MUX_WDOUT_sle<=0;
						MemWrite<=0;
						CMPsle<=0;
						ifj<=0;
						kuo<=0;
						start<=0;
						MULTsle<=0;
						M<=0;
						cp<=0;
						eret<=1;
						WA<=0;
					end
				endcase
			end
			
			6'b000001:begin
				case(IR[20:16])
					5'b00000:begin
						EXTsle<=0;
						npcsle<=1;
						MUX_ALU_B_sle<=0;
						ALUsle<=0;
						RegWrite<=0;
						Branch<=1;
						MUX_A3_sle<=0;
						MUX_WDOUT_sle<=0;
						MemWrite<=0;
						CMPsle<=5;
						ifj<=0;
						kuo<=0;
						start<=0;
						MULTsle<=0;
						M<=0;
						cp<=0;
						eret<=0;
						WA<=0;
					end/////bltz
					
					5'b00001:begin
						EXTsle<=0;
						npcsle<=1;
						MUX_ALU_B_sle<=0;
						ALUsle<=0;
						RegWrite<=0;
						Branch<=1;
						MUX_A3_sle<=0;
						MUX_WDOUT_sle<=0;
						MemWrite<=0;
						CMPsle<=2;
						ifj<=0;
						kuo<=0;
						start<=0;
						MULTsle<=0;
						M<=0;
						cp<=0;
						eret<=0;
						WA<=0;
					end/////bgez
					
					default begin
						EXTsle<=0;
						npcsle<=0;
						MUX_ALU_B_sle<=0;
						ALUsle<=0;
						RegWrite<=0;
						Branch<=0;
						MUX_A3_sle<=0;
						MUX_WDOUT_sle<=0;
						MemWrite<=0;
						CMPsle<=0;
						ifj<=0;
						kuo<=0;
						start<=0;
						MULTsle<=0;
						M<=0;
						cp<=0;
						eret<=0;
						WA<=0;
					end
				endcase
			end
			
					
			default begin
				EXTsle<=0;
				npcsle<=0;
				MUX_ALU_B_sle<=0;
				ALUsle<=0;
				RegWrite<=0;
				Branch<=0;
				MUX_A3_sle<=0;
				MUX_WDOUT_sle<=0;
				MemWrite<=0;
				CMPsle<=0;
				ifj<=0;
				kuo<=0;
				start<=0;
				MULTsle<=0;
				M<=0;
				cp<=0;
				eret<=0;
				WA<=1;
			end
		endcase
	end


endmodule
